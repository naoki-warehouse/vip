module main

struct IPv4Hdr {

}